/* Akshay Trikha
   MicroPs Lab 7
   November 6th, 2019
*/

/////////////////////////////////////////////
// aes
//   Top level module with SPI interface and SPI core
/////////////////////////////////////////////

module aes(input  logic clk,
           input  logic sck,
           input  logic sdi,
           output logic sdo,
           input  logic load,
           output logic done);

    logic [127:0] key, plainText, cypherText;

    aes_spi spi(sck, sdi, sdo, done, key, plainText, cypherText);
    aes_core core(clk, load, key, plainText, done, cypherText);
endmodule

/////////////////////////////////////////////
// aes_spi
//   SPI interface.  Shifts in key and plaintext
//   Captures cyphertext when done, then shifts it out
//   Tricky cases to properly change sdo on negedge clk
/////////////////////////////////////////////

module aes_spi(input  logic sck,
               input  logic sdi,
               output logic sdo,
               input  logic done,
               output logic [127:0] key, plainText,
               input  logic [127:0] cypherText);

    logic         sdodelayed, wasdone;
    logic [127:0] cyphertextcaptured;

    // assert load
    // apply 256 sclks to shift in key and plaintext, starting with plaintext[0]
    // then deassert load, wait until done
    // then apply 128 sclks to shift out cyphertext, starting with cyphertext[0]
    always_ff @(posedge sck)
        if (!wasdone)  {cyphertextcaptured, plainText, key} = {cypherText, plainText[126:0], key, sdi};
        else           {cyphertextcaptured, plainText, key} = {cyphertextcaptured[126:0], plainText, key, sdi};

    // sdo should change on the negative edge of sck
    always_ff @(negedge sck) begin
        wasdone = done;
        sdodelayed = cyphertextcaptured[126];
    end

    // when done is first asserted, shift out msb before clock edge
    assign sdo = (done & !wasdone) ? cypherText[127] : sdodelayed;
endmodule

/////////////////////////////////////////////
// aes_core
//   top level AES encryption module
//   when load is asserted, takes the current key and plaintext
//   generates cyphertext and asserts done when complete 11 cycles later
//
//   See FIPS-197 with Nk = 4, Nb = 4, Nr = 10
//
//   The key and message are 128-bit values packed into an array of 16 bytes as
//   shown below
//        [127:120] [95:88] [63:56] [31:24]     S0,0    S0,1    S0,2    S0,3
//        [119:112] [87:80] [55:48] [23:16]     S1,0    S1,1    S1,2    S1,3
//        [111:104] [79:72] [47:40] [15:8]      S2,0    S2,1    S2,2    S2,3
//        [103:96]  [71:64] [39:32] [7:0]       S3,0    S3,1    S3,2    S3,3
//
//   Equivalently, the values are packed into four words as given
//        [127:96]  [95:64] [63:32] [31:0]      w[0]    w[1]    w[2]    w[3]
/////////////////////////////////////////////

module aes_core(input  logic         clk,
                input  logic         load,
                input  logic [127:0] key,
                input  logic [127:0] plainText,
                output logic         done,
                output logic [127:0] cypherText);

      // internal logic for enable signals in control path
      logic cypherTextOn;
      logic subByteOn;
      logic shiftRowsOn;
      logic mixColumnsOn;
      logic keyExpansionOn;
      logic addRoundKeyOn;
		logic [3:0]currentRound; // current round #

      // internal logic for subByte and mux
      logic [127:0]noSubByte;
      logic [127:0]subByte;

      // internal logic for shiftRows and mux
      logic [127:0]noShiftRows;
      logic [127:0]shiftRows;

      // internal logic for mixColumns and mux
      logic [127:0]noMixColumns;
      logic [127:0]mixColumns;

      // internal logic for addRoundKey and mux
      logic [127:0]noAddRoundKey;
      logic [127:0]addRoundKey;

      // internal logic for keyExpansion and mux
      logic [127:0]oldKey;
      logic [127:0]newKey;
      logic [127:0]calculatedKey;

      // internal logic for done round flop
      logic [127:0]oldCypherText;

      // instantiating submodules
      controller    c1(clk, load, cypherTextOn, subByteOn, shiftRowsOn, mixColumnsOn, keyExpansionOn, addRoundKeyOn, currentRound, done);
      assign noSubByte = cypherTextOn ? plainText : cypherText;

      // use subByte transformation if subByteOn == 1
      subByte       sb1(noSubByte, subByte);
      assign noShiftRows = subByteOn ? subByte : noSubByte;

      // use shiftRows transformation if shiftRowsOn == 1
      shiftRows     sr1(noShiftRows, shiftRows);
      assign noMixColumns = shiftRowsOn ? shiftRows : noShiftRows;

      // use mixColumns transformation if mixColumnsOn == 1
      mixColumns    mc1(noMixColumns, mixColumns);
      assign noAddRoundKey = mixColumnsOn ? mixColumns : noMixColumns;

      // keyExpansion
      keyExpansion  k1(calculatedKey, currentRound, oldKey);
      assign calculatedKey = keyExpansionOn ? newKey : key;

      // use addRoundKey transformation if addRoundKeyOn == 1
      addRoundKey ar1(noAddRoundKey, calculatedKey, addRoundKey);
      assign oldCypherText = addRoundKeyOn ? addRoundKey : noAddRoundKey;
		// flip flop between oldKey and newKey on rising clock edge
	   always_ff @(posedge clk)
				newKey <= oldKey;

      // flip flop between oldCypherText and cypherText on rising clock edge
	   always_ff @(posedge clk)
				cypherText <= oldCypherText;

endmodule
